

* File includes subcircuits and technology definitions
.include ./SRAM_bits.cir


*this cell emulates load from SRAM cells,
* Number refers to the load from than number of cells
.subckt memLoad ttt fff number=254
Xnt ttt gnd dead nn ww='number*5'
Xnf fff gnd dead nn ww='number*5'
.ends memLoad




*********begin: topLevel*****

* Parameters
.global gnd vdd
.param gnd=0


*********begin: topLevel*****
.param per = 8ns
.param dataLead=500ps
.param lw=1358
.param wirew=12

vdd vdd 0 'supply'

Xclok clk               dat1 period='per' start='per+dataLead' total=1 duty=0.5 sz=50
Xrdwr rdw               dat1 period='per' start='2*per'        total=2 duty=1
Xdii din                dat1 period='per' start='per'          total=4 duty=2   sz=30



*Tied clk to din on dec model so that cho will be asserted
Xde1 cho clk clk decModel
Xwr1 bt1 bf1 din rdw clk write1
Xwi1 bt1 btt bf1 bff     wire_dual len='lw' wid='wirew'
Xml1 btt bff             memLoad number =31
Xme1 btt bff cho         mem1
Xsu1 btt bff set rst rdw clk readSub
*In the line below im doing some hand waving because normally I would want to
*have 8 write lines going into the read collect 8, however, I'm just demonstrating
*the worst case of a single furthest away mem cell
Xrc dot set rst vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd readcollect8

.ic V(la:tt)=0 V(la:ff)=1
.ic V(bt2)=1
.tran 1p 'per*10'






