* This file contains all the subcircuits to be used in SRAM256.cir

***** long channel VTP = -0.9, VTN = 0.8 *****
*.include modelcard/1um.pm
*.param supply = 5
*.param ll = 1u

****** 50nm models***


.include C:\Users\steph\OneDrive - Oregon State University\ECE 471\transistor_models\50nm.pm
.param supply =1

.param lambda=25nm
.param ll='2*lambda'

****** 16nm low power models***
*.include ./modelcard/PTM_LP/16nm.pm
*.param supply =0.9
*.param ll=16nm

****** 16nm high peformance models***
*.include ./modelcard/PTM_HP/16nm.pm
*.param supply =0.7
*.param ll=16nm


.subckt wire iot iof len=10 wid=10
.param rr=0.8
.param cc = '200e-15'
rt iot iof 'rr*len*50/(wid)'
cf iof  0  'cc*len*wid*50/1e6'

.ends

.subckt wire_dual lt rt lf rf len=10 wid=10
Xt lt rt wire len='len' wid='wid'
Xf lf rf wire len='len' wid='wid'
.ends

.subckt nn d g s  ww=100
mnfet d g s 0 nmos L=ll w='ww*ll'
.ends

.subckt pp d g s   ww=100
mpfet d g s vdd pmos L=ll w='ww*ll'
.ends


.subckt inv out inn size=30 beta=2
XPP out inn vdd pp ww='size*beta/(beta+1)'
XNN out inn gnd nn ww='size/(beta+1)'
.ends

.subckt nnd2 out in1 in0 size=30 beta=2
Xap0 out in0 vdd pp ww='beta*size/(beta+2)'
Xap1 out in1 vdd pp ww='beta*size/(beta+2)'
Xan0 out in0 nng nn ww='2*size/(beta+2)'
Xan1 nng in1 0   nn ww='2*size/(beta+2)'
.ends nnd2

.subckt nor2 out in1 in0 size=30 beta=2
Xap0 ppi in0 vdd pp ww='2*beta*size/(2*beta+1)'
Xap1 out in1 ppi pp ww='2*beta*size/(2*beta+1)'
Xan0 out in0 0 nn ww='1*size/(2*beta+1)'
Xan1 out in1 0   nn ww='1*size/(2*beta+1)'
.ends nor2

.subckt latch out inn clk clb size=15 beta=2
Xn inn clk qin nn ww='5'
Xp inn clb qin pp ww='10'

Xfp qin ggg vdd pp ww='5'
Xfn qin ggg gnd nn ww='5'

Xi ggg qin     inv size='size'
Xo out ggg     inv size='3*size'
.ends latch

.subckt flop qqq ddd clk
Xinve clb clk inv
Xflip int ddd clb clk latch
Xflop qqq int clk clb latch
.ends flop

.subckt reg8 ot7 ot6 ot5 ot4 ot3 ot2 ot1 ot0 in7 in6 in5 in4 in3 in2 in1 in0 clk
x7 ot7 in7 clk flop
x6 ot6 in6 clk flop
x5 ot5 in5 clk flop
x4 ot4 in4 clk flop
x3 ot3 in3 clk flop
x2 ot2 in2 clk flop
x1 ot1 in1 clk flop
x0 ot0 in0 clk flop
.ends reg8

.subckt dat1 out period=1ns start=1ns sz=50 total=5 duty=3
V0 j0  0  PULSE('supply' 0 'start' 10p 10p 'duty*period-10ps' 'total*period')
x7 out j0 inv size='sz'
.ends dat1

*generates different data stream on all eight channels, buffered output
.subckt dat8 o7 o6 o5 o4 o3 o2 o1 o0 per=1ns start=1ns size=50
V0 j0  0  PULSE(0 'supply' 'start' 10p 10p '0.5*per-10ps' 'per')
V1 j1  0  PULSE(0 'supply' 'start' 10p 10p '0.5*per-10ps' '2*per')
V2 j2  0  PULSE(0 'supply' 'start' 10p 10p '0.5*per-10ps' '3*per')
V3 j3  0  PULSE(0 'supply' 'start' 10p 10p '0.5*per-10ps' '4*per')
V4 j4  0  PULSE('supply' 0 'start' 10p 10p '0.5*per-10ps' '1*per')
V5 j5  0  PULSE('supply' 0 'start' 10p 10p '1*per-10ps' '2*per')
V6 j6  0  PULSE('supply' 0 'start' 10p 10p '1.5*per-10ps' '3*per')
V7 j7  0  PULSE('supply' 0 'start' 10p 10p '2*per-10ps' '4*per')
xb o7 o6 o5 o4 o3 o2 o1 o0 j7 j6 j5 j4 j3 j2 j1 j0 buf8 sz='size'
.ends dat8

.subckt buf8 ot7 ot6 ot5 ot4 ot3 ot2 ot1 ot0 in7 in6 in5 in4 in3 in2 in1 in0 sz=100
x7 ot7 in7 inv size='sz'
x6 ot6 in6 inv size='sz'
x5 ot5 in5 inv size='sz'
x4 ot4 in4 inv size='sz'
x3 ot3 in3 inv size='sz'
x2 ot2 in2 inv size='sz'
x1 ot1 in1 inv size='sz'
x0 ot0 in0 inv size='sz'
.ends buf8


.subckt nnd3 out in2 in1 in0 size=20 beta=2
Xp0 out in0 vdd pp ww='beta*size/(beta+3)'
Xp1 out in1 vdd pp ww='beta*size/(beta+3)'
Xp2 out in2 vdd pp ww='beta*size/(beta+3)'
Xn0 out in0 nn0 nn ww='3*size/(beta+3)'
Xn1 nn0 in1 nn1 nn ww='3*size/(beta+3)'
Xn2 nn1 in2 gnd nn ww='3*size/(beta+3)'
.ends

.subckt senseAmp ot1 ot0 in1 in0 eva size=40
Xn0 ot0 in0 ot1 eva nnd3 size ='size'
Xn1 ot1 in1 ot0 eva nnd3 size ='size'
.ends senseAmp

.subckt decModel cho din clk size=100 beta=2
Xin1 nn1 din 	 inv
Xpt2 nn2 nn1 vdd nnd2
Xdu2 dd1 nn1 gnd nnd2
Xpt3 nn3 nn2 gnd nor2
Xdu3 dd2 nn2 vdd nor2 size='3*size'
Xpt4 nn4 nn3 vdd nnd2
Xdu4 dd3 nn3 gnd nnd2 size='15*size'
*Xin5 nn5 nn4 	 inv
*commented out above inv because it buffered my input to be behind the example waveform
Xpt5 nn5 nn4 clk nnd2
Xin6 cho nn5 	 inv
.ends decModel
**ope off on dec model

.subckt decModel_v2 cho din clk size=100 beta=2
Xin1 nn1 din 	 inv
Xpt2 nn2 nn1 vdd nnd2
Xdu2 dd1 nn1 gnd nnd2
Xin2 nn3 nn2 	 inv
Xpt3 nn4 nn3 vdd nnd2
Xin3 nn5 nn4 	 inv
Xdu3 dd2 nn3 vdd nor2 size='3*size'
Xpt4 nn6 nn5 vdd nnd2
Xdu4 dd3 nn5 gnd nnd2 size='15*size'
*Xpt3 nn3 nn2 gnd nor2
*Xdu3 dd2 nn2 vdd nor2 size='3*size'
*Xpt4 nn4 nn3 vdd nnd2
*Xdu4 dd3 nn3 gnd nnd2 size='15*size'
*Xin5 nn5 nn4 	 inv
Xpt5 nn7 nn6 clk nnd2
Xin6 cho nn7 	 inv
.ends decModel_v2

.subckt write1 btt bff dit rwt clk size=30 beta=2
Xin1 nn1 rwt     inv
Xnd2 nn2 nn1 clk nnd2
Xin2 nn3 nn2     inv
Xnn2 nn4 nn3 gnd nn
Xnn3 btt dit nn4 nn
Xin3 nn5 dit     inv
Xnn4 bff nn5 nn4 nn
Xpp4 btt clk vdd pp
Xpp5 bff clk vdd pp
.ends write1

*try 1
*.subckt read1 btt bff dot rdw clk size=100 beta=2
*Xnd1 nn1 rdw clk nnd2
*Xin1 tri nn1     inv
*Xnd2 set tri btt res nnd3
*Xnd3 res tri bff set nnd3
*Xin3 nn2 set     inv
*Xin4 nn4 res     inv
*Xin5 nn3 nn2     inv
*Xpp5 nn5 nn3 vdd pp
*Xnn6 nn5 nn4 gnd nn
*Xin7 dot nn5 	 inv
*Xin6 nn5 dot 	 inv
*.ends read1

.subckt read1 btt bff dot rwt clk size=10
Xnd1 nn1 rwt clk nnd2 size='size'
Xin1 nn2 nn1     inv  size='size'
Xse1 fal tru bff btt  nn2 senseAmp size='5*size'
Xin2 nn3 fal     inv  size='2*size'
Xin3 nn4 nn3     inv  size='2*size'
Xin4 nn5 tru     inv  size='2*size'
Xpp5 nn6 nn4 vdd pp   ww='2*size'
Xnn5 gnd nn5 nn6 nn   ww='size'
Xin5 nn6 dot     inv  size='size'
Xin6 dot nn6     inv  size='2*size'
.ends read1

*adjusting width seems to force btt and bff down to gnd & vdd harder
*this makes sense due to current being directly proportional to width
*sized for beta=2
*sized with 5 from reference nn and pp transistors
.subckt mem1 btt bff ope wid=5
Xnn1 btt ope nn1 nn ww='wid'
Xnn2 bff ope nn2 nn ww='wid'
Xpp3 vdd nn2 nn1 pp ww='2*wid'
Xnn3 nn1 nn2 gnd nn ww='wid'
Xpp4 vdd nn1 nn2 pp ww='2*wid'
Xnn4 nn2 nn1 gnd nn ww='wid'
.end mem1

*read sub is dut (seems like changing sizes doesnt do anything to output)
*sized according to reference sense amp provided
.subckt readSub btt bff set rst rdw clk size=40 beta=2
Xnd1 nn1 rdw clk nnd2     size = 'size'
Xin1 tri nn1     inv  	  size = 'size'
*Xsa1 set rst btt bff trg senseAmp size = '20'
Xnd3 set tri btt rst nnd3 size='size'
Xnd4 rst tri bff set nnd3 size='size'
.ends readSub

.subckt readcollect8 nnn st7 rs7 st6 rs6 st5 rs5 st4 rs4 st3 rs3 st2 rs2 st1 rs1 st0 rs0 size=30 beta=2
Xnd7 aa7 st7 st6 nnd2
Xnd6 aa6 st5 st4 nnd2
Xnd5 aa5 st3 st2 nnd2
Xnd4 aa4 st1 st0 nnd2
Xin7 hi7 aa7     inv
Xin6 hi6 aa6     inv
Xin5 hi5 aa5     inv
Xin4 hi4 aa4 	 inv
Xpp7 dot hi7 vdd pp ww='2*size'
Xpp6 dot hi6 vdd pp ww='2*size'
Xpp5 dot hi5 vdd pp ww='2*size'
Xpp4 dot hi4 vdd pp ww='2*size'
Xnd3 io3 rs7 rs6 nnd2
Xnd2 io2 rs5 rs4 nnd2
Xnd1 io1 rs3 rs2 nnd2
Xnd0 io0 rs1 rs0 nnd2
Xnn3 dot io3 gnd nn
Xnn2 dot io2 gnd nn
Xnn1 dot io1 gnd nn
Xnn0 dot io0 gnd nn
*output state holder
Xinx dot nnn  	 inv
Xiny nnn dot     inv
.ends readcollect8

.subckt decode2 o11 o10 o01 o00 di1 di0 df1 df0

.ends


.subckt decode_nor16

.ends

.subckt decode_nnd16

.ends


.subckt decode_16and1

.ends decode_16and1


.subckt dmux256 o255 o223 0012 o001 dt7 dt6 dt5 d4 dt3 dt1 dt0

.ends dmux256






